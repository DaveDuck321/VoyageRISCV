module fence(
    input wire clk,

    output wire error
);

assign error = 1'b0;

// TODO

endmodule
